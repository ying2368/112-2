library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity lab13_G06 is
    Port ( clk : in std_logic;
           hex0 : out std_logic_vector(6 downto 0);
           hex1 : out std_logic_vector(6 downto 0);
           hex2 : out std_logic_vector(7 downto 0);
           hex3 : out std_logic_vector(6 downto 0));
end lab13_G06;

architecture Behavioral of lab13_G06 is
    signal minutes : integer range 0 to 59 := 59;
    signal seconds : integer range 0 to 59 := 57;
    signal clk_div : integer := 0;

    function seven_segment(input : integer) return std_logic_vector is
    begin
        case input is
            when 0 => return "1000000";
            when 1 => return "1111001";
            when 2 => return "0100100";
            when 3 => return "0110000";
            when 4 => return "0011001";
            when 5 => return "0010010";
            when 6 => return "0000010"; 
            when 7 => return "1111000"; 
            when 8 => return "0000000";
            when 9 => return "0010000";
            when others => return "1111111";
        end case;
    end function;

begin
    process(clk)
    begin
        if rising_edge(clk) then
            clk_div <= clk_div + 1;
            if clk_div = 50000000 then
                clk_div <= 0;
                if seconds = 59 then
                    seconds <= 0;
                    if minutes = 59 then
                        minutes <= 0;
                    else
                        minutes <= minutes + 1;
                    end if;
                else
                    seconds <= seconds + 1;
                end if;
            end if;
        end if;
    end process;

    hex0 <= seven_segment(seconds mod 10);
    hex1 <= seven_segment(seconds / 10);
    hex2 <= '0' & seven_segment(minutes mod 10);
    hex3 <= seven_segment(minutes / 10);

end Behavioral;
