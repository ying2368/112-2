library verilog;
use verilog.vl_types.all;
entity s1111442_lab08_2 is
    port(
        clk             : in     vl_logic;
        clrn            : in     vl_logic;
        Q               : out    vl_logic_vector(1 downto 0)
    );
end s1111442_lab08_2;
